`include "ethernet_frame_pkg.sv"
`include "axi_master_model.sv"
`include "AXI_interface.sv"
`include "rtl_struct.sv"
`include "eth_core.sv"
`include "eth_tx.sv"
`include "dma_controller_tx.sv"
//`include "AXI_master.sv"
`include "AXI_slave.sv"
`include "dma_fifo.sv"
